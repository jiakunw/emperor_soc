// emperor_i2c_pkg.sv

`ifndef EMPEROR_I2C_PKG
    `define EMPEROR_I2C_PKG

    `include "uvm_macros.svh"

    package emperor_i2c_pkg;
        import uvm_pkg::*;
    endpackage
`endif