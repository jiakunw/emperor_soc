// emperor_axi_lite_types.sv

`ifndef EMPEROR_AXI_LITE_TYPES
    `define EMPEROR_AXI_LITE_TYPES

    `include "uvm_macros.svh"
    `include "emperor_axi_lite_if.sv"

    package emperor_axi_lite_types;
        import uvm_pkg::*;
    endpackage
`endif